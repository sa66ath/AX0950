CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 120 30 100 9
0 74 1153 502
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
30 C:\Program Files\CM60S\BOM.DAT
0 7
0 74 1153 502
144179219 0
0
6 Title:
5 Name:
0
0
0
24
7 Ground~
168 746 306 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
10 Capacitor~
219 643 416 0 2 5
0 2 8
0
0 0 848 90
4 47uF
10 0 38 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
10 FW Bridge~
219 535 415 0 4 9
0 2 9 8 10
0
0 0 848 90
6 BRIDGE
32 -40 74 -32
2 D2
46 -50 60 -42
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
88 0 0 256 1 0 0 0
1 D
3618 0 0
0
0
7 Op Amp~
219 354 391 0 3 7
0 5 11 6
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
11 Signal Gen~
195 192 392 0 64 64
0 12 5 2 86 -8 8 0 0 0
0 0 0 0 0 0 0 1116471296 0 1101004800
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
0 70 0 20 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -20/20V
-25 -30 24 -22
2 V2
-7 -40 7 -32
0
0
30 %D %1 %2 DC 0 SIN(0 20 70 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
11 Signal Gen~
195 185 226 0 64 64
0 17 13 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1086953882
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
1 50 0 6.3 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -6.3/6.3V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 6.3 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
7 Op Amp~
219 347 225 0 3 7
0 13 16 15
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U2
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
6 Diode~
219 405 226 0 2 5
0 15 3
0
0 0 848 0
6 1N4007
-21 -18 21 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 1 0 0
1 D
3747 0 0
0
0
6 Diode~
219 408 303 0 2 5
0 2 15
0
0 0 848 512
6 1N4007
-21 -18 21 -10
2 D5
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 1 0 0
1 D
3549 0 0
0
0
10 Capacitor~
219 439 243 0 2 5
0 13 3
0
0 0 848 90
6 1000uF
3 0 45 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
10 Capacitor~
219 439 281 0 2 5
0 2 13
0
0 0 848 90
6 1000uF
1 0 43 8
2 C5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
9 I Source~
198 745 259 0 2 5
0 14 2
0
0 0 17264 0
4 100m
16 0 44 8
3 Is1
20 -10 41 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
8903 0 0
0
0
12 Zener Diode~
219 634 279 0 2 5
0 2 7
0
0 0 848 90
5 1N759
15 -2 50 6
2 D8
26 -12 40 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
100 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
12 NPN Trans:B~
219 636 234 0 3 7
0 3 7 14
0
0 0 848 90
3 NPN
-13 -26 8 -18
2 Q2
-9 -36 5 -28
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3363 0 0
0
0
10 Capacitor~
219 699 262 0 2 5
0 2 14
0
0 0 848 90
4 10uF
7 0 35 8
2 C6
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7668 0 0
0
0
9 Resistor~
219 378 461 0 2 5
0 5 4
0
0 0 880 90
3 100
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 378 410 0 2 5
0 4 6
0
0 0 880 90
3 100
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 424 478 0 2 5
0 5 9
0
0 0 880 0
4 2.2k
-15 -14 13 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 420 391 0 2 5
0 6 10
0
0 0 880 0
4 2.2k
-15 -14 13 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 355 341 0 2 5
0 11 6
0
0 0 880 0
7 1.4142k
-24 -14 25 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 300 387 0 2 5
0 12 11
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 293 221 0 2 5
0 17 16
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 348 175 0 2 5
0 16 15
0
0 0 880 0
7 1.4142k
-24 -14 25 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 580 259 0 2 5
0 7 3
0
0 0 880 180
3 470
-11 -14 10 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
37
1 0 2 0 0 4096 0 1 0 0 3 2
746 300
745 298
2 0 3 0 0 8192 0 24 0 0 27 3
562 259
546 259
546 224
0 0 2 0 0 8192 0 0 0 23 10 3
745 298
630 298
630 447
0 0 4 0 0 4224 0 0 0 5 0 7
378 434
499 434
499 470
501 470
501 438
539 438
539 446
1 2 4 0 0 0 0 17 16 0 0 2
378 428
378 443
1 0 5 0 0 4096 0 16 0 0 8 2
378 479
378 478
2 0 6 0 0 4096 0 17 0 0 14 2
378 392
380 391
0 1 5 0 0 8320 0 0 18 15 0 3
261 397
261 478
406 478
2 1 7 0 0 8320 0 13 24 0 0 3
634 269
634 259
598 259
1 1 2 0 0 0 0 3 2 0 0 4
537 443
537 447
643 447
643 425
3 2 8 0 0 8320 0 3 2 0 0 4
537 379
537 375
643 375
643 407
2 2 9 0 0 8320 0 3 18 0 0 4
505 411
449 411
449 478
442 478
2 4 10 0 0 12416 0 19 3 0 0 6
438 391
501 391
501 362
577 362
577 411
569 411
1 0 6 0 0 4096 0 19 0 0 16 2
402 391
380 391
2 1 5 0 0 0 0 5 4 0 0 2
223 397
336 397
2 3 6 0 0 8320 0 20 4 0 0 4
373 341
380 341
380 391
372 391
1 0 11 0 0 8320 0 20 0 0 18 3
337 341
321 341
321 387
2 2 11 0 0 0 0 4 21 0 0 4
336 385
326 385
326 387
318 387
1 1 12 0 0 4224 0 21 5 0 0 2
282 387
223 387
0 0 13 0 0 8320 0 0 0 33 30 3
242 231
242 262
439 262
1 0 2 0 0 0 0 15 0 0 23 4
699 271
699 293
700 293
700 298
2 0 14 0 0 4096 0 15 0 0 24 2
699 253
699 227
2 0 2 0 0 0 0 12 0 0 26 4
745 280
745 298
634 298
634 303
3 1 14 0 0 4224 0 14 12 0 0 3
652 227
745 227
745 238
2 2 7 0 0 0 0 13 14 0 0 2
634 269
634 250
0 1 2 0 0 4224 0 0 13 29 0 3
439 303
634 303
634 289
1 0 3 0 0 12416 0 14 0 0 31 7
616 227
603 227
603 224
435 224
435 231
435 231
435 226
2 0 15 0 0 8320 0 9 0 0 32 3
398 303
378 303
378 226
1 1 2 0 0 0 0 11 9 0 0 3
439 290
439 303
418 303
1 2 13 0 0 0 0 10 11 0 0 2
439 252
439 272
2 2 3 0 0 0 0 8 10 0 0 3
415 226
439 226
439 234
1 0 15 0 0 0 0 8 0 0 34 4
395 226
378 226
378 224
373 224
2 1 13 0 0 0 0 6 7 0 0 2
216 231
329 231
2 3 15 0 0 0 0 23 7 0 0 4
366 175
373 175
373 225
365 225
1 0 16 0 0 8320 0 23 0 0 36 3
330 175
314 175
314 221
2 2 16 0 0 0 0 7 22 0 0 4
329 219
319 219
319 221
311 221
1 1 17 0 0 4224 0 22 6 0 0 2
275 221
216 221
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1 0.001 0.0002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4130610 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
736 459
0 0 0 0 0 0
12401 0
4 1 1
1
580 259
0 0 0 0 0	24 0 0 0
3213132 8550464 100 100 0 0
77 66 1127 336
0 502 1153 930
1127 66
77 66
1127 66
1127 336
740 298
1 0 0.054 0 1 1
12401 0
4 0.3 2e+016
1
580 259
0 0 0 0 0	24 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
