CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
28 104 1124 900
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
30 C:\Program Files\CM60S\BOM.DAT
0 7
28 104 1124 900
144179219 0
0
6 Title:
5 Name:
0
0
0
4
7 Ground~
168 553 515 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
9 V Source~
197 507 446 0 2 5
0 4 2
0
0 0 17264 0
3 280
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
4441 0 0
0
0
9 I Source~
198 603 453 0 2 5
0 3 2
0
0 0 17264 0
5 1.7mA
13 0 48 8
3 Is1
20 -10 41 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
3618 0 0
0
0
9 Resistor~
219 604 391 0 2 5
0 3 4
0
0 0 880 90
3 47k
4 0 25 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
4
1 0 2 0 0 4096 0 1 0 0 2 2
553 509
553 478
2 2 2 0 0 8320 0 3 2 0 0 4
603 474
603 478
507 478
507 467
1 1 3 0 0 4224 0 4 3 0 0 4
604 409
604 424
603 424
603 432
1 2 4 0 0 8320 0 2 4 0 0 4
507 425
507 365
604 365
604 373
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3540062 1210432 100 100 0 0
0 0 0 0
1 72 162 142
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 100 300
1
604 391
0 0 0 0 0	4 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
