CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 190 30 100 9
0 74 1157 557
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
30 C:\Program Files\CM60S\BOM.DAT
0 7
0 74 1157 557
144179219 0
0
6 Title:
5 Name:
0
0
0
12
6 Diode~
219 476 312 0 2 5
0 3 4
0
0 0 848 180
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 1 0 0
1 D
8953 0 0
0
0
7 Op Amp~
219 317 312 0 3 7
0 2 8 7
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 0 0 0 0
1 U
4441 0 0
0
0
7 Ground~
168 680 448 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 634 362 0 2 5
0 2 5
0
0 0 848 90
4 10uF
8 0 36 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 513 367 0 2 5
0 2 3
0
0 0 848 90
4 10uF
8 0 36 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
11 Signal Gen~
195 144 312 0 19 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1135869952
20
1 50 0 360 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -360/360V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 360 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
9 Resistor~
219 321 264 0 2 5
0 8 7
0
0 0 880 0
5 141.5
-17 -14 18 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 259 308 0 2 5
0 9 8
0
0 0 880 0
3 100
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 682 396 0 3 5
0 2 6 -1
0
0 0 880 90
3 10k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 679 342 0 2 5
0 6 5
0
0 0 880 90
3 47k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 587 311 0 2 5
0 3 5
0
0 0 880 0
3 15k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 419 311 0 2 5
0 7 4
0
0 0 880 0
4 220k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
16
2 0 3 0 0 4096 0 5 0 0 3 2
513 358
513 312
2 2 4 0 0 4224 0 12 1 0 0 4
437 311
458 311
458 312
466 312
1 1 3 0 0 4224 0 1 11 0 0 4
486 312
561 312
561 311
569 311
1 0 2 0 0 4096 0 4 0 0 8 2
634 371
634 425
2 0 5 0 0 4096 0 4 0 0 11 2
634 353
634 311
0 2 2 0 0 8192 0 0 6 7 0 3
291 380
291 317
175 317
0 1 2 0 0 8320 0 0 2 8 0 5
515 425
515 380
291 380
291 318
299 318
0 1 2 0 0 0 0 0 5 9 0 3
682 425
513 425
513 376
1 1 2 0 0 0 0 9 3 0 0 4
682 414
682 434
680 434
680 442
2 1 6 0 0 4224 0 9 10 0 0 4
682 378
682 368
679 368
679 360
2 2 5 0 0 8320 0 10 11 0 0 3
679 324
679 311
605 311
1 0 7 0 0 4224 0 12 0 0 13 3
401 311
346 311
346 312
3 2 7 0 0 0 0 2 7 0 0 4
335 312
347 312
347 264
339 264
2 1 8 0 0 8320 0 2 7 0 0 4
299 306
295 306
295 264
303 264
2 2 8 0 0 0 0 8 2 0 0 4
277 308
291 308
291 306
299 306
1 1 9 0 0 4224 0 6 8 0 0 4
175 307
233 307
233 308
241 308
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2230188 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 0.1
1
657 311
0 5 0 0 2	0 11 0 0
2623304 8550464 100 100 0 0
77 66 1127 336
0 502 1157 930
1127 66
77 66
1127 66
1127 336
0 0
10 0 -7.10543e-015 -54 10 10
12401 0
4 0.03 10000
1
500 312
0 3 0 0 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
