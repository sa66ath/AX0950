CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 200 30 100 9
138 315 1334 684
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
138 315 1334 684
144179219 0
0
6 Title:
5 Name:
0
0
0
34
11 Signal Gen~
195 39 404 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1008981771
20
1 1000 0 0.01 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -10m/10mV
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 10m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
10 Capacitor~
219 565 320 0 2 5
0 6 7
0
0 0 848 90
2 5n
12 0 26 8
2 C8
12 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
10 Capacitor~
219 615 299 0 2 5
0 6 5
0
0 0 848 0
4 500p
-14 -18 14 -10
2 C7
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Capacitor~
219 403 292 0 2 5
0 7 10
0
0 0 848 180
3 22n
-11 -18 10 -10
2 C6
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 403 351 0 2 5
0 9 8
0
0 0 848 180
3 22n
-11 -18 10 -10
2 C5
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
7 Ground~
168 1021 248 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 863 244 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 478 262 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
10 Capacitor~
219 864 209 0 2 5
0 2 12
0
0 0 848 90
4 50uF
8 0 36 8
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
10 Capacitor~
219 478 235 0 2 5
0 2 17
0
0 0 848 90
4 50uF
8 0 36 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
10 Capacitor~
219 402 444 0 2 5
0 2 16
0
0 0 848 90
4 330u
8 0 36 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
10 Capacitor~
219 203 444 0 2 5
0 2 15
0
0 0 848 90
4 680n
8 0 36 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
7 Ground~
168 95 516 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3834 0 0
0
0
9 V Source~
197 1019 192 0 2 5
0 12 2
0
0 0 17264 0
4 265V
10 0 38 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3363 0 0
0
0
7 Triode~
219 787 384 0 3 7
0 12 13 11
0
0 0 848 0
5 12AX7
23 0 58 8
3 V2B
30 -10 51 -2
0
0
14 %D %1 %2 %3 %S
0
0
4 VT-9
10

0 6 7 8 1 2 3 6 7 8
0
88 0 0 0 2 2 2 0
1 V
7668 0 0
0
0
7 Triode~
219 690 383 0 3 7
0 13 5 14
0
0 0 848 0
5 12AX7
23 0 58 8
3 V2A
30 -10 51 -2
0
0
14 %D %1 %2 %3 %S
0
0
4 VT-9
10

0 1 2 3 1 2 3 6 7 8
0
88 0 0 0 2 1 2 0
1 V
4718 0 0
0
0
7 Triode~
219 350 387 0 3 7
0 8 2 16
0
0 0 848 0
5 12AX7
23 0 58 8
3 V1B
30 -10 51 -2
0
0
14 %D %1 %2 %3 %S
0
0
4 VT-9
10

0 6 7 8 1 2 3 6 7 8
0
88 0 0 0 2 2 1 0
1 V
3874 0 0
0
0
7 Triode~
219 173 386 0 3 7
0 10 4 15
0
0 0 848 0
5 12AX7
23 0 58 8
3 V1A
30 -10 51 -2
0
0
14 %D %1 %2 %3 %S
0
0
4 VT-9
10

0 1 2 3 1 2 3 6 7 8
393221
88 0 0 0 2 1 1 0
1 V
6671 0 0
0
0
9 Resistor~
219 616 358 0 2 5
0 5 6
0
0 0 880 180
3 47k
-11 -14 10 -6
3 R15
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 621 438 0 2 5
0 5 3
0
0 0 880 180
3 47k
-11 -14 10 -6
3 R14
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 527 324 0 2 5
0 6 7
0
0 0 880 90
1 1
13 0 20 8
3 R13
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 527 404 0 3 5
0 2 6 -1
0
0 0 880 90
4 1meg
4 0 32 8
3 R12
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 474 414 0 2 5
0 3 9
0
0 0 880 90
4 1meg
4 0 32 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 474 463 0 3 5
0 2 3 -1
0
0 0 880 90
1 1
14 0 21 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 689 320 0 2 5
0 13 12
0
0 0 880 90
4 100k
1 0 29 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 566 163 0 2 5
0 12 17
0
0 0 880 180
3 10k
-11 -14 10 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 352 263 0 2 5
0 8 17
0
0 0 880 90
4 100k
1 0 29 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 171 265 0 2 5
0 10 17
0
0 0 880 90
4 100k
1 0 29 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 349 445 0 3 5
0 2 16 -1
0
0 0 880 90
3 820
5 0 26 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 777 445 0 3 5
0 2 11 -1
0
0 0 880 90
4 100k
1 0 29 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 678 446 0 3 5
0 2 14 -1
0
0 0 880 90
3 820
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 306 441 0 3 5
0 2 2 -1
0
0 0 880 90
2 1M
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 162 444 0 3 5
0 2 15 -1
0
0 0 880 90
4 2700
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 92 441 0 3 5
0 2 4 -1
0
0 0 880 90
2 1M
8 0 22 8
3 R16
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
49
0 0 2 0 0 12288 0 0 0 35 33 4
306 387
306 419
269 419
269 502
2 1 3 0 0 4224 0 20 23 0 0 3
603 438
474 438
474 432
2 1 2 0 0 0 0 1 34 0 0 5
70 409
83 409
83 467
92 467
92 459
0 1 4 0 0 4096 0 0 1 45 0 2
92 399
70 399
2 1 5 0 0 8320 0 3 19 0 0 4
624 299
642 299
642 358
634 358
1 0 6 0 0 8320 0 3 0 0 9 3
606 299
586 299
586 358
1 0 6 0 0 0 0 2 0 0 9 4
565 329
565 354
527 354
527 359
0 2 7 0 0 8192 0 0 2 18 0 4
525 292
525 301
565 301
565 311
2 0 6 0 0 144 0 19 0 0 17 4
598 358
542 358
542 359
527 359
1 2 5 0 0 0 0 19 16 0 0 4
634 358
656 358
656 383
664 383
1 2 5 0 0 128 0 20 16 0 0 4
639 438
656 438
656 383
664 383
2 0 8 0 0 4096 0 5 0 0 48 2
394 351
352 351
1 0 2 0 0 0 0 24 0 0 27 2
474 481
474 497
1 2 3 0 0 128 0 23 24 0 0 2
474 432
474 445
1 2 9 0 0 4224 0 5 23 0 0 3
412 351
474 351
474 396
1 0 2 0 0 0 0 22 0 0 27 2
527 422
527 497
1 2 6 0 0 0 0 21 22 0 0 2
527 342
527 386
1 2 7 0 0 4224 0 4 21 0 0 3
412 292
527 292
527 306
2 0 10 0 0 4224 0 4 0 0 49 2
394 292
173 292
1 0 2 0 0 8192 0 30 0 0 27 3
777 463
777 496
678 496
3 2 11 0 0 4224 0 15 30 0 0 4
776 407
776 419
777 419
777 427
1 0 12 0 0 4096 0 15 0 0 43 2
787 358
787 163
0 2 13 0 0 4224 0 0 15 25 0 4
690 350
753 350
753 384
761 384
2 0 12 0 0 0 0 25 0 0 43 2
689 302
689 163
1 1 13 0 0 0 0 16 25 0 0 4
690 357
690 346
689 346
689 338
3 2 14 0 0 4224 0 16 31 0 0 4
679 406
679 420
678 420
678 428
1 0 2 0 0 8192 0 31 0 0 33 4
678 464
678 497
395 497
395 502
1 0 2 0 0 0 0 12 0 0 33 2
203 453
203 502
2 0 15 0 0 8320 0 12 0 0 46 3
203 435
203 422
162 422
1 0 2 0 0 0 0 33 0 0 33 2
162 462
162 502
1 0 2 0 0 0 0 32 0 0 33 4
306 459
306 497
307 497
307 502
1 0 2 0 0 0 0 29 0 0 33 4
349 463
349 497
350 497
350 502
1 1 2 0 0 8320 0 11 13 0 0 4
402 453
402 502
95 502
95 510
2 0 16 0 0 8320 0 11 0 0 47 3
402 435
402 418
349 418
2 2 2 0 0 128 0 17 32 0 0 3
324 387
306 387
306 423
2 0 17 0 0 8320 0 28 0 0 37 4
171 247
171 162
352 162
352 163
0 2 17 0 0 0 0 0 27 42 0 3
478 163
352 163
352 245
1 1 2 0 0 0 0 10 8 0 0 2
478 244
478 256
1 1 2 0 0 0 0 9 7 0 0 4
864 218
864 230
863 230
863 238
2 1 2 0 0 0 0 14 6 0 0 4
1019 213
1019 234
1021 234
1021 242
2 0 12 0 0 0 0 9 0 0 43 2
864 200
864 163
2 2 17 0 0 0 0 10 26 0 0 3
478 226
478 163
548 163
1 1 12 0 0 4224 0 26 14 0 0 3
584 163
1019 163
1019 171
1 1 2 0 0 0 0 34 13 0 0 4
92 459
92 502
95 502
95 510
2 2 4 0 0 8320 0 34 18 0 0 3
92 423
92 386
147 386
3 2 15 0 0 0 0 18 33 0 0 2
162 409
162 426
2 3 16 0 0 0 0 29 17 0 0 4
349 427
349 418
339 418
339 410
1 1 8 0 0 4224 0 27 17 0 0 4
352 281
352 353
350 353
350 361
1 1 10 0 0 0 0 18 28 0 0 4
173 360
173 291
171 291
171 283
0
0
25 0 1
0
0
0
0 0 0
0
0 0 0
40 1 20 20000
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
3605162 1210432 100 100 0 0
77 66 1169 276
139 313 300 383
1169 66
77 66
1169 66
1169 276
0 0
20000 20 5 4.46189e+270 19980 30
12401 0
4 1 200
1
777 429
0 11 0 0 2	30 0 0 0
3802020 8550464 100 100 0 0
77 66 1157 276
138 684 1334 1053
1157 66
77 66
1157 66
1157 276
0 0
0.005 0 0.24 -0.24 0.005 0.005
12401 0
4 1e-006 5
1
655 358
0 5 0 0 1	0 10 0 0
528238 4683840 100 100 0 0
77 66 1169 276
138 684 1332 1053
592 66
1169 66
1169 78
1169 110
0 0
519.835 20000 -43.1429 -52.5714 19980 19980
12403 0
4 5000 30
1
352 338
0 8 0 0 1	0 48 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
