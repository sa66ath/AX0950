CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 210 30 100 9
0 74 1157 502
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
30 C:\Program Files\CM60S\BOM.DAT
0 7
0 74 1157 502
144179219 0
0
6 Title:
5 Name:
0
0
0
15
10 Capacitor~
219 498 398 0 2 5
0 2 4
0
0 0 848 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
10 Capacitor~
219 569 396 0 2 5
0 2 3
0
0 0 848 90
4 10uF
8 0 36 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
7 Ground~
168 565 486 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
6 Diode~
219 385 396 0 2 5
0 6 5
0
0 0 848 692
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 1 0 0
1 D
6153 0 0
0
0
7 Op Amp~
219 316 437 0 3 7
0 2 8 6
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U2
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
5394 0 0
0
0
6 Diode~
219 385 312 0 2 5
0 7 5
0
0 0 848 692
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 1 0 0
1 D
7734 0 0
0
0
7 Op Amp~
219 320 311 0 3 7
0 2 9 7
0
0 0 848 0
5 IDEAL
-21 -31 14 -23
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
11 Signal Gen~
195 144 312 0 19 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1135869952
20
1 50 0 360 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -360/360V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 360 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
9 Resistor~
219 522 348 0 2 5
0 4 3
0
0 0 880 0
4 1Meg
-13 -14 15 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 472 349 0 2 5
0 5 4
0
0 0 880 0
4 1Meg
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 643 379 0 3 5
0 2 3 -1
0
0 0 880 90
4 220k
2 0 30 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 335 397 0 2 5
0 8 6
0
0 0 880 0
3 100
-10 -14 11 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 267 431 0 2 5
0 7 8
0
0 0 880 0
3 100
-10 -14 11 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 321 264 0 2 5
0 9 7
0
0 0 880 0
5 141.5
-17 -14 18 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 259 308 0 2 5
0 10 9
0
0 0 880 0
3 100
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
25
0 2 3 0 0 4224 0 0 11 13 0 3
565 352
643 352
643 361
2 0 3 0 0 0 0 9 0 0 13 2
540 348
565 349
1 0 2 0 0 4096 0 1 0 0 6 2
498 407
498 458
2 0 4 0 0 4224 0 1 0 0 5 2
498 389
498 348
1 2 4 0 0 0 0 9 10 0 0 4
504 348
498 348
498 349
490 349
0 0 2 0 0 8192 0 0 0 0 12 4
434 411
434 458
522 458
522 463
0 0 5 0 0 4096 0 0 0 0 8 2
434 393
434 349
1 0 5 0 0 4096 0 10 0 0 14 4
454 349
408 349
408 350
403 350
1 0 2 0 0 4096 0 5 0 0 20 2
298 443
197 443
1 2 2 0 0 4096 0 7 8 0 0 2
302 317
175 317
1 1 2 0 0 0 0 11 3 0 0 4
643 397
643 472
565 472
565 480
1 1 2 0 0 0 0 2 3 0 0 6
569 405
569 463
522 463
522 463
565 463
565 480
2 0 3 0 0 0 0 2 0 0 0 4
569 387
569 364
565 364
565 349
2 2 5 0 0 8320 0 6 4 0 0 4
395 312
403 312
403 396
395 396
1 2 6 0 0 4096 0 4 12 0 0 4
375 396
361 396
361 397
353 397
1 0 7 0 0 12416 0 13 0 0 21 5
249 431
245 431
245 346
348 346
348 311
3 2 6 0 0 8320 0 5 12 0 0 4
334 437
347 437
347 397
353 397
2 1 8 0 0 8320 0 5 12 0 0 4
298 431
295 431
295 397
317 397
2 2 8 0 0 0 0 13 5 0 0 2
285 431
298 431
1 2 2 0 0 8320 0 3 8 0 0 8
565 480
565 476
196 476
196 506
197 506
197 377
175 377
175 317
1 0 7 0 0 128 0 6 0 0 22 5
375 312
348 312
348 311
346 311
346 312
3 2 7 0 0 0 0 7 14 0 0 6
338 311
346 311
346 312
347 312
347 264
339 264
2 1 9 0 0 8320 0 7 14 0 0 4
302 305
295 305
295 264
303 264
2 2 9 0 0 0 0 15 7 0 0 4
277 308
291 308
291 305
302 305
1 1 10 0 0 4224 0 8 15 0 0 4
175 307
233 307
233 308
241 308
0
0
17 0 2
0
0
0
0 0 0
0
0 0 0
3 0 1 4
19 20 0.004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2557286 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 3 20
0
3343702 8550464 100 100 0 0
77 66 1127 336
0 502 1157 930
1127 66
77 66
1127 66
1127 336
0 0
20 19 0.00035 -7e-005 0.999994 0.999994
12401 0
4 3 2000
1
456 349
0 5 0 0 1	10 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
